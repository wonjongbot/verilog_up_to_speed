`default_nettype none

module thruwire( input logic i_sw,
                 output logic o_led);
    assign o_led = i_sw;
endmodule
